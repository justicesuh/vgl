module gl43

#flag  -I @VROOT/thirdparty/glad
#flag @VROOT/thirdparty/glad/glad.o
#include <glad.h>

import const (
	GL_ACTIVE_RESOURCES
	GL_ACTIVE_VARIABLES
	GL_ANY_SAMPLES_PASSED_CONSERVATIVE
	GL_ARRAY_SIZE
	GL_ARRAY_STRIDE
	GL_ATOMIC_COUNTER_BUFFER_INDEX
	GL_ATOMIC_COUNTER_BUFFER_REFERENCED_BY_COMPUTE_SHADER
	GL_AUTO_GENERATE_MIPMAP
	GL_BLOCK_INDEX
	GL_BUFFER
	GL_BUFFER_BINDING
	GL_BUFFER_DATA_SIZE
	GL_BUFFER_VARIABLE
	GL_CAVEAT_SUPPORT
	GL_CLEAR_BUFFER
	GL_COLOR_COMPONENTS
	GL_COLOR_ENCODING
	GL_COLOR_RENDERABLE
	GL_COMPRESSED_R11_EAC
	GL_COMPRESSED_RG11_EAC
	GL_COMPRESSED_RGB8_ETC2
	GL_COMPRESSED_RGB8_PUNCHTHROUGH_ALPHA1_ETC2
	GL_COMPRESSED_RGBA8_ETC2_EAC
	GL_COMPRESSED_SIGNED_R11_EAC
	GL_COMPRESSED_SIGNED_RG11_EAC
	GL_COMPRESSED_SRGB8_ALPHA8_ETC2_EAC
	GL_COMPRESSED_SRGB8_ETC2
	GL_COMPRESSED_SRGB8_PUNCHTHROUGH_ALPHA1_ETC2
	GL_COMPUTE_SHADER
	GL_COMPUTE_SHADER_BIT
	GL_COMPUTE_SUBROUTINE
	GL_COMPUTE_SUBROUTINE_UNIFORM
	GL_COMPUTE_TEXTURE
	GL_COMPUTE_WORK_GROUP_SIZE
	GL_CONTEXT_FLAG_DEBUG_BIT
	GL_DEBUG_CALLBACK_FUNCTION
	GL_DEBUG_CALLBACK_USER_PARAM
	GL_DEBUG_GROUP_STACK_DEPTH
	GL_DEBUG_LOGGED_MESSAGES
	GL_DEBUG_NEXT_LOGGED_MESSAGE_LENGTH
	GL_DEBUG_OUTPUT
	GL_DEBUG_OUTPUT_SYNCHRONOUS
	GL_DEBUG_SEVERITY_HIGH
	GL_DEBUG_SEVERITY_LOW
	GL_DEBUG_SEVERITY_MEDIUM
	GL_DEBUG_SEVERITY_NOTIFICATION
	GL_DEBUG_SOURCE_API
	GL_DEBUG_SOURCE_APPLICATION
	GL_DEBUG_SOURCE_OTHER
	GL_DEBUG_SOURCE_SHADER_COMPILER
	GL_DEBUG_SOURCE_THIRD_PARTY
	GL_DEBUG_SOURCE_WINDOW_SYSTEM
	GL_DEBUG_TYPE_DEPRECATED_BEHAVIOR
	GL_DEBUG_TYPE_ERROR
	GL_DEBUG_TYPE_MARKER
	GL_DEBUG_TYPE_OTHER
	GL_DEBUG_TYPE_PERFORMANCE
	GL_DEBUG_TYPE_POP_GROUP
	GL_DEBUG_TYPE_PORTABILITY
	GL_DEBUG_TYPE_PUSH_GROUP
	GL_DEBUG_TYPE_UNDEFINED_BEHAVIOR
	GL_DEPTH_COMPONENTS
	GL_DEPTH_RENDERABLE
	GL_DEPTH_STENCIL_TEXTURE_MODE
	GL_DISPATCH_INDIRECT_BUFFER
	GL_DISPATCH_INDIRECT_BUFFER_BINDING
	GL_DISPLAY_LIST
	GL_FILTER
	GL_FRAGMENT_SUBROUTINE
	GL_FRAGMENT_SUBROUTINE_UNIFORM
	GL_FRAGMENT_TEXTURE
	GL_FRAMEBUFFER_BLEND
	GL_FRAMEBUFFER_DEFAULT_FIXED_SAMPLE_LOCATIONS
	GL_FRAMEBUFFER_DEFAULT_HEIGHT
	GL_FRAMEBUFFER_DEFAULT_LAYERS
	GL_FRAMEBUFFER_DEFAULT_SAMPLES
	GL_FRAMEBUFFER_DEFAULT_WIDTH
	GL_FRAMEBUFFER_RENDERABLE
	GL_FRAMEBUFFER_RENDERABLE_LAYERED
	GL_FULL_SUPPORT
	GL_GEOMETRY_SUBROUTINE
	GL_GEOMETRY_SUBROUTINE_UNIFORM
	GL_GEOMETRY_TEXTURE
	GL_GET_TEXTURE_IMAGE_FORMAT
	GL_GET_TEXTURE_IMAGE_TYPE
	GL_IMAGE_CLASS_1_X_16
	GL_IMAGE_CLASS_1_X_32
	GL_IMAGE_CLASS_1_X_8
	GL_IMAGE_CLASS_10_10_10_2
	GL_IMAGE_CLASS_11_11_10
	GL_IMAGE_CLASS_2_X_16
	GL_IMAGE_CLASS_2_X_32
	GL_IMAGE_CLASS_2_X_8
	GL_IMAGE_CLASS_4_X_16
	GL_IMAGE_CLASS_4_X_32
	GL_IMAGE_CLASS_4_X_8
	GL_IMAGE_COMPATIBILITY_CLASS
	GL_IMAGE_PIXEL_FORMAT
	GL_IMAGE_PIXEL_TYPE
	GL_IMAGE_TEXEL_SIZE
	GL_INTERNALFORMAT_ALPHA_SIZE
	GL_INTERNALFORMAT_ALPHA_TYPE
	GL_INTERNALFORMAT_BLUE_SIZE
	GL_INTERNALFORMAT_BLUE_TYPE
	GL_INTERNALFORMAT_DEPTH_SIZE
	GL_INTERNALFORMAT_DEPTH_TYPE
	GL_INTERNALFORMAT_GREEN_SIZE
	GL_INTERNALFORMAT_GREEN_TYPE
	GL_INTERNALFORMAT_PREFERRED
	GL_INTERNALFORMAT_RED_SIZE
	GL_INTERNALFORMAT_RED_TYPE
	GL_INTERNALFORMAT_SHARED_SIZE
	GL_INTERNALFORMAT_STENCIL_SIZE
	GL_INTERNALFORMAT_STENCIL_TYPE
	GL_INTERNALFORMAT_SUPPORTED
	GL_IS_PER_PATCH
	GL_IS_ROW_MAJOR
	GL_LOCATION
	GL_LOCATION_INDEX
	GL_MANUAL_GENERATE_MIPMAP
	GL_MATRIX_STRIDE
	GL_MAX_COMBINED_COMPUTE_UNIFORM_COMPONENTS
	GL_MAX_COMBINED_DIMENSIONS
	GL_MAX_COMBINED_SHADER_OUTPUT_RESOURCES
	GL_MAX_COMBINED_SHADER_STORAGE_BLOCKS
	GL_MAX_COMPUTE_ATOMIC_COUNTER_BUFFERS
	GL_MAX_COMPUTE_ATOMIC_COUNTERS
	GL_MAX_COMPUTE_IMAGE_UNIFORMS
	GL_MAX_COMPUTE_SHADER_STORAGE_BLOCKS
	GL_MAX_COMPUTE_SHARED_MEMORY_SIZE
	GL_MAX_COMPUTE_TEXTURE_IMAGE_UNITS
	GL_MAX_COMPUTE_UNIFORM_BLOCKS
	GL_MAX_COMPUTE_UNIFORM_COMPONENTS
	GL_MAX_COMPUTE_WORK_GROUP_COUNT
	GL_MAX_COMPUTE_WORK_GROUP_INVOCATIONS
	GL_MAX_COMPUTE_WORK_GROUP_SIZE
	GL_MAX_DEBUG_GROUP_STACK_DEPTH
	GL_MAX_DEBUG_LOGGED_MESSAGES
	GL_MAX_DEBUG_MESSAGE_LENGTH
	GL_MAX_DEPTH
	GL_MAX_ELEMENT_INDEX
	GL_MAX_FRAGMENT_SHADER_STORAGE_BLOCKS
	GL_MAX_FRAMEBUFFER_HEIGHT
	GL_MAX_FRAMEBUFFER_LAYERS
	GL_MAX_FRAMEBUFFER_SAMPLES
	GL_MAX_FRAMEBUFFER_WIDTH
	GL_MAX_GEOMETRY_SHADER_STORAGE_BLOCKS
	GL_MAX_HEIGHT
	GL_MAX_LABEL_LENGTH
	GL_MAX_LAYERS
	GL_MAX_NAME_LENGTH
	GL_MAX_NUM_ACTIVE_VARIABLES
	GL_MAX_NUM_COMPATIBLE_SUBROUTINES
	GL_MAX_SHADER_STORAGE_BLOCK_SIZE
	GL_MAX_SHADER_STORAGE_BUFFER_BINDINGS
	GL_MAX_TESS_CONTROL_SHADER_STORAGE_BLOCKS
	GL_MAX_TESS_EVALUATION_SHADER_STORAGE_BLOCKS
	GL_MAX_UNIFORM_LOCATIONS
	GL_MAX_VERTEX_ATTRIB_BINDINGS
	GL_MAX_VERTEX_ATTRIB_RELATIVE_OFFSET
	GL_MAX_VERTEX_SHADER_STORAGE_BLOCKS
	GL_MAX_WIDTH
	GL_MIPMAP
	GL_NAME_LENGTH
	GL_NUM_ACTIVE_VARIABLES
	GL_NUM_SHADING_LANGUAGE_VERSIONS
	GL_OFFSET
	GL_PRIMITIVE_RESTART_FIXED_INDEX
	GL_PROGRAM
	GL_PROGRAM_INPUT
	GL_PROGRAM_OUTPUT
	GL_PROGRAM_PIPELINE
	GL_QUERY
	GL_READ_PIXELS
	GL_READ_PIXELS_FORMAT
	GL_READ_PIXELS_TYPE
	GL_REFERENCED_BY_COMPUTE_SHADER
	GL_REFERENCED_BY_FRAGMENT_SHADER
	GL_REFERENCED_BY_GEOMETRY_SHADER
	GL_REFERENCED_BY_TESS_CONTROL_SHADER
	GL_REFERENCED_BY_TESS_EVALUATION_SHADER
	GL_REFERENCED_BY_VERTEX_SHADER
	GL_SAMPLER
	GL_SHADER
	GL_SHADER_IMAGE_ATOMIC
	GL_SHADER_IMAGE_LOAD
	GL_SHADER_IMAGE_STORE
	GL_SHADER_STORAGE_BARRIER_BIT
	GL_SHADER_STORAGE_BLOCK
	GL_SHADER_STORAGE_BUFFER
	GL_SHADER_STORAGE_BUFFER_BINDING
	GL_SHADER_STORAGE_BUFFER_OFFSET_ALIGNMENT
	GL_SHADER_STORAGE_BUFFER_SIZE
	GL_SHADER_STORAGE_BUFFER_START
	GL_SIMULTANEOUS_TEXTURE_AND_DEPTH_TEST
	GL_SIMULTANEOUS_TEXTURE_AND_DEPTH_WRITE
	GL_SIMULTANEOUS_TEXTURE_AND_STENCIL_TEST
	GL_SIMULTANEOUS_TEXTURE_AND_STENCIL_WRITE
	GL_SRGB_READ
	GL_SRGB_WRITE
	GL_STENCIL_COMPONENTS
	GL_STENCIL_RENDERABLE
	GL_TESS_CONTROL_SUBROUTINE
	GL_TESS_CONTROL_SUBROUTINE_UNIFORM
	GL_TESS_CONTROL_TEXTURE
	GL_TESS_EVALUATION_SUBROUTINE
	GL_TESS_EVALUATION_SUBROUTINE_UNIFORM
	GL_TESS_EVALUATION_TEXTURE
	GL_TEXTURE_BUFFER_OFFSET
	GL_TEXTURE_BUFFER_OFFSET_ALIGNMENT
	GL_TEXTURE_BUFFER_SIZE
	GL_TEXTURE_COMPRESSED_BLOCK_HEIGHT
	GL_TEXTURE_COMPRESSED_BLOCK_SIZE
	GL_TEXTURE_COMPRESSED_BLOCK_WIDTH
	GL_TEXTURE_GATHER
	GL_TEXTURE_GATHER_SHADOW
	GL_TEXTURE_IMAGE_FORMAT
	GL_TEXTURE_IMAGE_TYPE
	GL_TEXTURE_IMMUTABLE_LEVELS
	GL_TEXTURE_SHADOW
	GL_TEXTURE_VIEW
	GL_TEXTURE_VIEW_MIN_LAYER
	GL_TEXTURE_VIEW_MIN_LEVEL
	GL_TEXTURE_VIEW_NUM_LAYERS
	GL_TEXTURE_VIEW_NUM_LEVELS
	GL_TOP_LEVEL_ARRAY_SIZE
	GL_TOP_LEVEL_ARRAY_STRIDE
	GL_TRANSFORM_FEEDBACK_VARYING
	GL_TYPE
	GL_UNIFORM
	GL_UNIFORM_BLOCK
	GL_UNIFORM_BLOCK_REFERENCED_BY_COMPUTE_SHADER
	GL_VERTEX_ATTRIB_ARRAY_LONG
	GL_VERTEX_ATTRIB_BINDING
	GL_VERTEX_ATTRIB_RELATIVE_OFFSET
	GL_VERTEX_BINDING_BUFFER
	GL_VERTEX_BINDING_DIVISOR
	GL_VERTEX_BINDING_OFFSET
	GL_VERTEX_BINDING_STRIDE
	GL_VERTEX_SUBROUTINE
	GL_VERTEX_SUBROUTINE_UNIFORM
	GL_VERTEX_TEXTURE
	GL_VIEW_CLASS_128_BITS
	GL_VIEW_CLASS_16_BITS
	GL_VIEW_CLASS_24_BITS
	GL_VIEW_CLASS_32_BITS
	GL_VIEW_CLASS_48_BITS
	GL_VIEW_CLASS_64_BITS
	GL_VIEW_CLASS_8_BITS
	GL_VIEW_CLASS_96_BITS
	GL_VIEW_CLASS_BPTC_FLOAT
	GL_VIEW_CLASS_BPTC_UNORM
	GL_VIEW_CLASS_RGTC1_RED
	GL_VIEW_CLASS_RGTC2_RG
	GL_VIEW_CLASS_S3TC_DXT1_RGB
	GL_VIEW_CLASS_S3TC_DXT1_RGBA
	GL_VIEW_CLASS_S3TC_DXT3_RGBA
	GL_VIEW_CLASS_S3TC_DXT5_RGBA
	GL_VIEW_COMPATIBILITY_CLASS
)

pub fn bind_vertex_buffer(bindingindex int, buffer int, offset i64, stride int) {
	C.glBindVertexBuffer(bindingindex, buffer, offset, stride)
}

pub fn clear_buffer_data(target int, internalformat int, format int, type int, data []f32) {
	C.glClearBufferData(target, internalformat, format, type, data)
}

pub fn clear_buffer_data(target int, internalformat int, format int, type int, data []int) {
	C.glClearBufferData(target, internalformat, format, type, data)
}

pub fn clear_buffer_data(target int, internalformat int, format int, type int, data []i16) {
	C.glClearBufferData(target, internalformat, format, type, data)
}

pub fn clear_buffer_data(target int, internalformat int, format int, type int, data voidptr) {
	C.glClearBufferData(target, internalformat, format, type, data)
}

pub fn clear_buffer_data(target int, internalformat int, format int, type int, data voidptr) {
	C.glClearBufferData(target, internalformat, format, type, data)
}

pub fn clear_buffer_data(target int, internalformat int, format int, type int, data voidptr) {
	C.glClearBufferData(target, internalformat, format, type, data)
}

pub fn clear_buffer_data(target int, internalformat int, format int, type int, data voidptr) {
	C.glClearBufferData(target, internalformat, format, type, data)
}

pub fn clear_buffer_sub_data(target int, internalformat int, offset i64, size i64, format int, type int, data []f32) {
	C.glClearBufferSubData(target, internalformat, offset, size, format, type, data)
}

pub fn clear_buffer_sub_data(target int, internalformat int, offset i64, size i64, format int, type int, data []int) {
	C.glClearBufferSubData(target, internalformat, offset, size, format, type, data)
}

pub fn clear_buffer_sub_data(target int, internalformat int, offset i64, size i64, format int, type int, data []i16) {
	C.glClearBufferSubData(target, internalformat, offset, size, format, type, data)
}

pub fn clear_buffer_sub_data(target int, internalformat int, offset i64, size i64, format int, type int, data voidptr) {
	C.glClearBufferSubData(target, internalformat, offset, size, format, type, data)
}

pub fn clear_buffer_sub_data(target int, internalformat int, offset i64, size i64, format int, type int, data voidptr) {
	C.glClearBufferSubData(target, internalformat, offset, size, format, type, data)
}

pub fn clear_buffer_sub_data(target int, internalformat int, offset i64, size i64, format int, type int, data voidptr) {
	C.glClearBufferSubData(target, internalformat, offset, size, format, type, data)
}

pub fn clear_buffer_sub_data(target int, internalformat int, offset i64, size i64, format int, type int, data voidptr) {
	C.glClearBufferSubData(target, internalformat, offset, size, format, type, data)
}

pub fn copy_image_sub_data(src_name int, src_target int, src_level int, src_x int, src_y int, src_z int, dst_name int, dst_target int, dst_level int, dst_x int, dst_y int, dst_z int, src_width int, src_height int, src_depth int) {
	C.glCopyImageSubData(src_name, src_target, src_level, src_x, src_y, src_z, dst_name, dst_target, dst_level, dst_x, dst_y, dst_z, src_width, src_height, src_depth)
}

pub fn debug_message_callback(